** sch_path: /home/gaston/Documents/simulacion.sch
.subckt simulacion

V1 net1 GND 1.8
V2 in GND PULSE(0 1.8 0 1n 1n 5n 10n 4)
R1 out GND 1k m=1
x1 net1 in out GND inversor
**** begin user architecture code
.lib /home/gaston/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt



.control
tran 0.5n 40n
write std_not4_tb.raw
.endc
.save all


**** end user architecture code
.ends

* expanding   symbol:  /home/gaston/Documents/inversor.sym # of pins=4
** sym_path: /home/gaston/Documents/inversor.sym
** sch_path: /home/gaston/Documents/inversor.sch
.subckt inversor Vdd Vin Vout Vss
*.PININFO Vdd:I Vss:I Vin:I Vout:O
XM2 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2.1 nf=1 m=1
XM1 Vout Vin Vss Vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.05 nf=1 m=1
.ends

.GLOBAL GND
